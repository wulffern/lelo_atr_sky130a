magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect 0 0 3328 2560
use LELOATR_NCH_12CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1664 480
use LELOATR_NCH_12C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1664 1280
use LELOATR_NCH_12C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1664 2080
use LELOATR_NCH_12CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1664 2560
use LELOATR_NCH_12CTAPBOT xb1 
transform 1 0 1664 0 1 0
box 1664 0 3328 480
use LELOATR_NCH_12C1F2 xb2 
transform 1 0 1664 0 1 480
box 1664 480 3328 1280
use LELOATR_NCH_12C5F0 xb3 
transform 1 0 1664 0 1 1280
box 1664 1280 3328 2080
use LELOATR_NCH_12CTAPTOP xb4 
transform 1 0 1664 0 1 2080
box 1664 2080 3328 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 3328 2560
<< end >>
