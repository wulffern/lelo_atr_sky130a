magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1848 928
<< pdiff >>
rect 416 200 1248 280
rect 416 280 1248 360
rect 416 360 1248 440
rect 416 440 1248 520
rect 416 520 1248 600
<< ptap >>
rect -96 -40 96 40
rect 1568 -40 1760 40
rect -96 40 96 120
rect 1568 40 1760 120
rect -96 120 96 200
rect 1568 120 1760 200
rect -96 200 96 280
rect 1568 200 1760 280
rect -96 280 96 360
rect 1568 280 1760 360
rect -96 360 96 440
rect 1568 360 1760 440
rect -96 440 96 520
rect 1568 440 1760 520
rect -96 520 96 600
rect 1568 520 1760 600
rect -96 600 96 680
rect 1568 600 1760 680
rect -96 680 96 760
rect 1568 680 1760 760
rect -96 760 96 840
rect 1568 760 1760 840
<< poly >>
rect 160 -22 1504 22
rect 160 138 1504 182
rect 160 298 1504 342
rect 160 458 1504 502
rect 160 618 1504 662
rect 160 778 1504 822
rect 160 280 224 360
rect 1440 280 1504 360
rect 160 360 224 440
rect 1440 360 1504 440
rect 160 440 224 520
rect 1440 440 1504 520
<< m1 >>
rect 160 360 224 440
rect 288 600 480 680
rect 1184 40 1376 120
rect 160 40 224 120
rect 288 40 480 120
rect 1184 40 1376 120
rect 160 120 224 200
rect 288 120 480 200
rect 1184 120 1376 200
rect 160 200 224 280
rect 288 200 480 280
rect 1184 200 1376 280
rect 160 280 224 360
rect 288 280 480 360
rect 1184 280 1376 360
rect 160 360 224 440
rect 288 360 480 440
rect 1184 360 1376 440
rect 160 440 224 520
rect 288 440 480 520
rect 1184 440 1376 520
rect 160 520 224 600
rect 288 520 480 600
rect 1184 520 1376 600
rect 160 600 224 680
rect 288 600 480 680
rect 1184 600 1376 680
rect 160 680 224 760
rect 288 680 480 760
rect 1184 680 1376 760
<< pcontact >>
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 1451 300 1493 320
rect 1451 320 1493 340
rect 1451 340 1493 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 1451 360 1493 380
rect 1451 380 1493 400
rect 1451 400 1493 420
rect 1451 420 1493 440
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 1451 440 1493 460
rect 1451 460 1493 480
rect 1451 480 1493 500
<< locali >>
rect -96 -40 96 40
rect 1568 -40 1760 40
rect -96 40 96 120
rect 1568 40 1760 120
rect -96 120 96 200
rect 1568 120 1760 200
rect -96 200 96 280
rect 288 200 1248 280
rect 1568 200 1760 280
rect -96 280 96 360
rect 160 280 224 360
rect 1440 280 1504 360
rect 1568 280 1760 360
rect -96 360 96 440
rect -96 360 96 440
rect 160 360 224 440
rect 416 360 1376 440
rect 1440 360 1504 440
rect 1568 360 1760 440
rect -96 440 96 520
rect 160 440 224 520
rect 1440 440 1504 520
rect 1568 440 1760 520
rect -96 520 96 600
rect 288 520 1248 600
rect 1568 520 1760 600
rect -96 600 96 680
rect 1568 600 1760 680
rect -96 680 96 760
rect 1568 680 1760 760
rect -96 760 96 840
rect 1568 760 1760 840
<< ptapc >>
rect -32 200 32 280
rect 1632 200 1696 280
rect -32 280 32 360
rect 1632 280 1696 360
rect -32 360 32 440
rect 1632 360 1696 440
rect -32 440 32 520
rect 1632 440 1696 520
rect -32 520 32 600
rect 1632 520 1696 600
<< ndcontact >>
rect 448 220 480 240
rect 448 240 480 260
rect 480 220 544 240
rect 480 240 544 260
rect 544 220 608 240
rect 544 240 608 260
rect 608 220 672 240
rect 608 240 672 260
rect 672 220 736 240
rect 672 240 736 260
rect 736 220 800 240
rect 736 240 800 260
rect 800 220 864 240
rect 800 240 864 260
rect 864 220 928 240
rect 864 240 928 260
rect 928 220 992 240
rect 928 240 992 260
rect 992 220 1056 240
rect 992 240 1056 260
rect 1056 220 1120 240
rect 1056 240 1120 260
rect 1120 220 1184 240
rect 1120 240 1184 260
rect 1184 220 1216 240
rect 1184 240 1216 260
rect 448 380 480 400
rect 448 400 480 420
rect 480 380 544 400
rect 480 400 544 420
rect 544 380 608 400
rect 544 400 608 420
rect 608 380 672 400
rect 608 400 672 420
rect 672 380 736 400
rect 672 400 736 420
rect 736 380 800 400
rect 736 400 800 420
rect 800 380 864 400
rect 800 400 864 420
rect 864 380 928 400
rect 864 400 928 420
rect 928 380 992 400
rect 928 400 992 420
rect 992 380 1056 400
rect 992 400 1056 420
rect 1056 380 1120 400
rect 1056 400 1120 420
rect 1120 380 1184 400
rect 1120 400 1184 420
rect 1184 380 1216 400
rect 1184 400 1216 420
rect 448 540 480 560
rect 448 560 480 580
rect 480 540 544 560
rect 480 560 544 580
rect 544 540 608 560
rect 544 560 608 580
rect 608 540 672 560
rect 608 560 672 580
rect 672 540 736 560
rect 672 560 736 580
rect 736 540 800 560
rect 736 560 800 580
rect 800 540 864 560
rect 800 560 864 580
rect 864 540 928 560
rect 864 560 928 580
rect 928 540 992 560
rect 928 560 992 580
rect 992 540 1056 560
rect 992 560 1056 580
rect 1056 540 1120 560
rect 1056 560 1120 580
rect 1120 540 1184 560
rect 1120 560 1184 580
rect 1184 540 1216 560
rect 1184 560 1216 580
<< viali >>
rect 320 208 352 216
rect 320 216 352 224
rect 320 224 352 232
rect 320 232 352 240
rect 320 240 352 248
rect 320 248 352 256
rect 320 256 352 264
rect 320 264 352 272
rect 352 208 416 216
rect 352 216 416 224
rect 352 224 416 232
rect 352 232 416 240
rect 352 240 416 248
rect 352 248 416 256
rect 352 256 416 264
rect 352 264 416 272
rect 416 208 448 216
rect 416 216 448 224
rect 416 224 448 232
rect 416 232 448 240
rect 416 240 448 248
rect 416 248 448 256
rect 416 256 448 264
rect 416 264 448 272
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 1216 368 1248 376
rect 1216 376 1248 384
rect 1216 384 1248 392
rect 1216 392 1248 400
rect 1216 400 1248 408
rect 1216 408 1248 416
rect 1216 416 1248 424
rect 1216 424 1248 432
rect 1248 368 1312 376
rect 1248 376 1312 384
rect 1248 384 1312 392
rect 1248 392 1312 400
rect 1248 400 1312 408
rect 1248 408 1312 416
rect 1248 416 1312 424
rect 1248 424 1312 432
rect 1312 368 1344 376
rect 1312 376 1344 384
rect 1312 384 1344 392
rect 1312 392 1344 400
rect 1312 400 1344 408
rect 1312 408 1344 416
rect 1312 416 1344 424
rect 1312 424 1344 432
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 320 528 352 536
rect 320 536 352 544
rect 320 544 352 552
rect 320 552 352 560
rect 320 560 352 568
rect 320 568 352 576
rect 320 576 352 584
rect 320 584 352 592
rect 352 528 416 536
rect 352 536 416 544
rect 352 544 416 552
rect 352 552 416 560
rect 352 560 416 568
rect 352 568 416 576
rect 352 576 416 584
rect 352 584 416 592
rect 416 528 448 536
rect 416 536 448 544
rect 416 544 448 552
rect 416 552 448 560
rect 416 560 448 568
rect 416 568 448 576
rect 416 576 448 584
rect 416 584 448 592
<< pwell >>
rect -184 -128 1848 928
<< labels >>
flabel m1 s 160 360 224 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 288 600 480 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -96 360 96 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 1184 40 1376 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -184 -128 1848 928
<< end >>
