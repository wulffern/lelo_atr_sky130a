magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect 0 0 2304 2560
use LELOATR_NCH_4CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1152 480
use LELOATR_NCH_4C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1152 1280
use LELOATR_NCH_4C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1152 2080
use LELOATR_NCH_4CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1152 2560
use LELOATR_NCH_4CTAPBOT xb1 
transform 1 0 1152 0 1 0
box 1152 0 2304 480
use LELOATR_NCH_4C1F2 xb2 
transform 1 0 1152 0 1 480
box 1152 480 2304 1280
use LELOATR_NCH_4C5F0 xb3 
transform 1 0 1152 0 1 1280
box 1152 1280 2304 2080
use LELOATR_NCH_4CTAPTOP xb4 
transform 1 0 1152 0 1 2080
box 1152 2080 2304 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 2304 2560
<< end >>
