magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1208 608
<< ntap >>
rect -96 120 1120 200
rect -96 200 1120 280
rect -96 280 1120 360
rect -96 360 96 440
rect 928 360 1120 440
rect -96 440 96 520
rect 928 440 1120 520
<< locali >>
rect -96 120 1120 200
rect -96 200 1120 280
rect -96 280 1120 360
rect -96 360 96 440
rect 928 360 1120 440
rect -96 440 96 520
rect 928 440 1120 520
<< ntapc >>
rect 160 200 800 280
<< nwell >>
rect -184 -128 1208 608
<< labels >>
<< properties >>
string FIXED_BBOX -184 -128 1208 608
<< end >>
