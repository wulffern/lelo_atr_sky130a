magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1208 928
<< pdiff >>
rect 416 200 608 280
rect 416 280 608 360
rect 416 360 608 440
rect 416 440 608 520
rect 416 520 608 600
<< ntap >>
rect -96 -40 96 40
rect 928 -40 1120 40
rect -96 40 96 120
rect 928 40 1120 120
rect -96 120 96 200
rect 928 120 1120 200
rect -96 200 96 280
rect 928 200 1120 280
rect -96 280 96 360
rect 928 280 1120 360
rect -96 360 96 440
rect 928 360 1120 440
rect -96 440 96 520
rect 928 440 1120 520
rect -96 520 96 600
rect 928 520 1120 600
rect -96 600 96 680
rect 928 600 1120 680
rect -96 680 96 760
rect 928 680 1120 760
rect -96 760 96 840
rect 928 760 1120 840
<< poly >>
rect 160 -22 864 22
rect 160 138 864 182
rect 160 298 864 342
rect 160 458 864 502
rect 160 618 864 662
rect 160 778 864 822
rect 160 280 224 360
rect 800 280 864 360
rect 160 360 224 440
rect 800 360 864 440
rect 160 440 224 520
rect 800 440 864 520
<< m1 >>
rect 160 360 224 440
rect 288 600 480 680
rect 544 40 736 120
rect 160 40 224 120
rect 288 40 480 120
rect 544 40 736 120
rect 160 120 224 200
rect 288 120 480 200
rect 544 120 736 200
rect 160 200 224 280
rect 288 200 480 280
rect 544 200 736 280
rect 160 280 224 360
rect 288 280 480 360
rect 544 280 736 360
rect 160 360 224 440
rect 288 360 480 440
rect 544 360 736 440
rect 160 440 224 520
rect 288 440 480 520
rect 544 440 736 520
rect 160 520 224 600
rect 288 520 480 600
rect 544 520 736 600
rect 160 600 224 680
rect 288 600 480 680
rect 544 600 736 680
rect 160 680 224 760
rect 288 680 480 760
rect 544 680 736 760
<< pcontact >>
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 811 300 853 320
rect 811 320 853 340
rect 811 340 853 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 811 360 853 380
rect 811 380 853 400
rect 811 400 853 420
rect 811 420 853 440
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 811 440 853 460
rect 811 460 853 480
rect 811 480 853 500
<< locali >>
rect -96 -40 96 40
rect 928 -40 1120 40
rect -96 40 96 120
rect 928 40 1120 120
rect -96 120 96 200
rect 928 120 1120 200
rect -96 200 96 280
rect 288 200 608 280
rect 928 200 1120 280
rect -96 280 96 360
rect 160 280 224 360
rect 800 280 864 360
rect 928 280 1120 360
rect -96 360 96 440
rect -96 360 96 440
rect 160 360 224 440
rect 416 360 736 440
rect 800 360 864 440
rect 928 360 1120 440
rect -96 440 96 520
rect 160 440 224 520
rect 800 440 864 520
rect 928 440 1120 520
rect -96 520 96 600
rect 288 520 608 600
rect 928 520 1120 600
rect -96 600 96 680
rect 928 600 1120 680
rect -96 680 96 760
rect 928 680 1120 760
rect -96 760 96 840
rect 928 760 1120 840
<< ntapc >>
rect -32 200 32 280
rect 992 200 1056 280
rect -32 280 32 360
rect 992 280 1056 360
rect -32 360 32 440
rect 992 360 1056 440
rect -32 440 32 520
rect 992 440 1056 520
rect -32 520 32 600
rect 992 520 1056 600
<< pdcontact >>
rect 448 220 480 240
rect 448 240 480 260
rect 480 220 544 240
rect 480 240 544 260
rect 544 220 576 240
rect 544 240 576 260
rect 448 380 480 400
rect 448 400 480 420
rect 480 380 544 400
rect 480 400 544 420
rect 544 380 576 400
rect 544 400 576 420
rect 448 540 480 560
rect 448 560 480 580
rect 480 540 544 560
rect 480 560 544 580
rect 544 540 576 560
rect 544 560 576 580
<< viali >>
rect 320 208 352 216
rect 320 216 352 224
rect 320 224 352 232
rect 320 232 352 240
rect 320 240 352 248
rect 320 248 352 256
rect 320 256 352 264
rect 320 264 352 272
rect 352 208 416 216
rect 352 216 416 224
rect 352 224 416 232
rect 352 232 416 240
rect 352 240 416 248
rect 352 248 416 256
rect 352 256 416 264
rect 352 264 416 272
rect 416 208 448 216
rect 416 216 448 224
rect 416 224 448 232
rect 416 232 448 240
rect 416 240 448 248
rect 416 248 448 256
rect 416 256 448 264
rect 416 264 448 272
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 576 368 608 376
rect 576 376 608 384
rect 576 384 608 392
rect 576 392 608 400
rect 576 400 608 408
rect 576 408 608 416
rect 576 416 608 424
rect 576 424 608 432
rect 608 368 672 376
rect 608 376 672 384
rect 608 384 672 392
rect 608 392 672 400
rect 608 400 672 408
rect 608 408 672 416
rect 608 416 672 424
rect 608 424 672 432
rect 672 368 704 376
rect 672 376 704 384
rect 672 384 704 392
rect 672 392 704 400
rect 672 400 704 408
rect 672 408 704 416
rect 672 416 704 424
rect 672 424 704 432
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 320 528 352 536
rect 320 536 352 544
rect 320 544 352 552
rect 320 552 352 560
rect 320 560 352 568
rect 320 568 352 576
rect 320 576 352 584
rect 320 584 352 592
rect 352 528 416 536
rect 352 536 416 544
rect 352 544 416 552
rect 352 552 416 560
rect 352 560 416 568
rect 352 568 416 576
rect 352 576 416 584
rect 352 584 416 592
rect 416 528 448 536
rect 416 536 448 544
rect 416 544 448 552
rect 416 552 448 560
rect 416 560 448 568
rect 416 568 448 576
rect 416 576 448 584
rect 416 584 448 592
<< nwell >>
rect -184 -128 1208 928
<< labels >>
flabel m1 s 160 360 224 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 288 600 480 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -96 360 96 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 544 40 736 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -184 -128 1208 928
<< end >>
