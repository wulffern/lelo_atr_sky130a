magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect 0 0 2816 2560
use LELOATR_PCH_8CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1408 480
use LELOATR_PCH_8C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1408 1280
use LELOATR_PCH_8C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1408 2080
use LELOATR_PCH_8CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1408 2560
use LELOATR_PCH_8CTAPBOT xb1 
transform 1 0 1408 0 1 0
box 1408 0 2816 480
use LELOATR_PCH_8C1F2 xb2 
transform 1 0 1408 0 1 480
box 1408 480 2816 1280
use LELOATR_PCH_8C5F0 xb3 
transform 1 0 1408 0 1 1280
box 1408 1280 2816 2080
use LELOATR_PCH_8CTAPTOP xb4 
transform 1 0 1408 0 1 2080
box 1408 2080 2816 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 2816 2560
<< end >>
