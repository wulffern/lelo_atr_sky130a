magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1208 608
<< ntap >>
rect -96 -40 96 40
rect 928 -40 1120 40
rect -96 40 96 120
rect 928 40 1120 120
rect -96 120 1120 200
rect -96 200 1120 280
rect -96 280 1120 360
<< locali >>
rect -96 -40 96 40
rect 928 -40 1120 40
rect -96 40 96 120
rect 928 40 1120 120
rect -96 120 1120 200
rect -96 200 1120 280
rect -96 280 1120 360
<< ntapc >>
rect 160 200 864 280
<< nwell >>
rect -184 -128 1208 608
<< labels >>
<< properties >>
string FIXED_BBOX -184 -128 1208 608
<< end >>
