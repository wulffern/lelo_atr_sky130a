magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1336 928
<< pdiff >>
rect 416 40 736 120
rect 416 120 736 200
rect 416 200 736 280
rect 416 280 736 360
rect 416 360 736 440
rect 416 440 736 520
rect 416 520 736 600
rect 416 600 736 680
rect 416 680 736 760
<< ntap >>
rect -96 -40 96 40
rect 1056 -40 1248 40
rect -96 40 96 120
rect 1056 40 1248 120
rect -96 120 96 200
rect 1056 120 1248 200
rect -96 200 96 280
rect 1056 200 1248 280
rect -96 280 96 360
rect 1056 280 1248 360
rect -96 360 96 440
rect 1056 360 1248 440
rect -96 440 96 520
rect 1056 440 1248 520
rect -96 520 96 600
rect 1056 520 1248 600
rect -96 600 96 680
rect 1056 600 1248 680
rect -96 680 96 760
rect 1056 680 1248 760
rect -96 760 96 840
rect 1056 760 1248 840
<< poly >>
rect 160 146 992 334
rect 160 466 992 654
rect 160 -22 992 22
rect 160 200 224 280
rect 928 200 992 280
rect 160 280 224 360
rect 928 280 992 360
rect 160 360 224 440
rect 928 360 992 440
rect 160 440 224 520
rect 928 440 992 520
rect 160 520 224 600
rect 928 520 992 600
rect 160 778 992 822
<< m1 >>
rect 160 360 224 440
rect 288 600 480 680
rect 672 40 864 120
rect 160 40 224 120
rect 288 40 480 120
rect 672 40 864 120
rect 160 120 224 200
rect 288 120 480 200
rect 672 120 864 200
rect 160 200 224 280
rect 288 200 480 280
rect 672 200 864 280
rect 160 280 224 360
rect 288 280 480 360
rect 672 280 864 360
rect 160 360 224 440
rect 288 360 480 440
rect 672 360 864 440
rect 160 440 224 520
rect 288 440 480 520
rect 672 440 864 520
rect 160 520 224 600
rect 288 520 480 600
rect 672 520 864 600
rect 160 600 224 680
rect 288 600 480 680
rect 672 600 864 680
rect 160 680 224 760
rect 288 680 480 760
rect 672 680 864 760
<< pcontact >>
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 939 300 981 320
rect 939 320 981 340
rect 939 340 981 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 939 360 981 380
rect 939 380 981 400
rect 939 400 981 420
rect 939 420 981 440
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 939 440 981 460
rect 939 460 981 480
rect 939 480 981 500
<< locali >>
rect -96 -40 96 40
rect 1056 -40 1248 40
rect -96 40 96 120
rect 288 40 736 120
rect 1056 40 1248 120
rect -96 120 96 200
rect 1056 120 1248 200
rect -96 200 96 280
rect 1056 200 1248 280
rect -96 280 96 360
rect 160 280 224 360
rect 928 280 992 360
rect 1056 280 1248 360
rect -96 360 96 440
rect -96 360 96 440
rect 160 360 224 440
rect 416 360 864 440
rect 928 360 992 440
rect 1056 360 1248 440
rect -96 440 96 520
rect 160 440 224 520
rect 928 440 992 520
rect 1056 440 1248 520
rect -96 520 96 600
rect 1056 520 1248 600
rect -96 600 96 680
rect 1056 600 1248 680
rect -96 680 96 760
rect 288 680 736 760
rect 1056 680 1248 760
rect -96 760 96 840
rect 1056 760 1248 840
<< ntapc >>
rect -32 200 32 280
rect 1120 200 1184 280
rect -32 280 32 360
rect 1120 280 1184 360
rect -32 360 32 440
rect 1120 360 1184 440
rect -32 440 32 520
rect 1120 440 1184 520
rect -32 520 32 600
rect 1120 520 1184 600
<< pdcontact >>
rect 448 60 480 80
rect 448 80 480 100
rect 480 60 544 80
rect 480 80 544 100
rect 544 60 608 80
rect 544 80 608 100
rect 608 60 672 80
rect 608 80 672 100
rect 672 60 704 80
rect 672 80 704 100
rect 448 380 480 400
rect 448 400 480 420
rect 480 380 544 400
rect 480 400 544 420
rect 544 380 608 400
rect 544 400 608 420
rect 608 380 672 400
rect 608 400 672 420
rect 672 380 704 400
rect 672 400 704 420
rect 448 700 480 720
rect 448 720 480 740
rect 480 700 544 720
rect 480 720 544 740
rect 544 700 608 720
rect 544 720 608 740
rect 608 700 672 720
rect 608 720 672 740
rect 672 700 704 720
rect 672 720 704 740
<< viali >>
rect 320 48 352 56
rect 320 56 352 64
rect 320 64 352 72
rect 320 72 352 80
rect 320 80 352 88
rect 320 88 352 96
rect 320 96 352 104
rect 320 104 352 112
rect 352 48 416 56
rect 352 56 416 64
rect 352 64 416 72
rect 352 72 416 80
rect 352 80 416 88
rect 352 88 416 96
rect 352 96 416 104
rect 352 104 416 112
rect 416 48 448 56
rect 416 56 448 64
rect 416 64 448 72
rect 416 72 448 80
rect 416 80 448 88
rect 416 88 448 96
rect 416 96 448 104
rect 416 104 448 112
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 704 368 736 376
rect 704 376 736 384
rect 704 384 736 392
rect 704 392 736 400
rect 704 400 736 408
rect 704 408 736 416
rect 704 416 736 424
rect 704 424 736 432
rect 736 368 800 376
rect 736 376 800 384
rect 736 384 800 392
rect 736 392 800 400
rect 736 400 800 408
rect 736 408 800 416
rect 736 416 800 424
rect 736 424 800 432
rect 800 368 832 376
rect 800 376 832 384
rect 800 384 832 392
rect 800 392 832 400
rect 800 400 832 408
rect 800 408 832 416
rect 800 416 832 424
rect 800 424 832 432
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 320 688 352 696
rect 320 696 352 704
rect 320 704 352 712
rect 320 712 352 720
rect 320 720 352 728
rect 320 728 352 736
rect 320 736 352 744
rect 320 744 352 752
rect 352 688 416 696
rect 352 696 416 704
rect 352 704 416 712
rect 352 712 416 720
rect 352 720 416 728
rect 352 728 416 736
rect 352 736 416 744
rect 352 744 416 752
rect 416 688 448 696
rect 416 696 448 704
rect 416 704 448 712
rect 416 712 448 720
rect 416 720 448 728
rect 416 728 448 736
rect 416 736 448 744
rect 416 744 448 752
<< pmoslvt >>
rect 416 146 736 334
rect 416 466 736 654
<< nwell >>
rect -184 -128 1336 928
<< labels >>
flabel m1 s 160 360 224 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 288 600 480 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -96 360 96 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 672 40 864 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -184 -128 1336 928
<< end >>
