magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1592 928
<< pdiff >>
rect 416 40 992 120
rect 416 120 992 200
rect 416 200 992 280
rect 416 280 992 360
rect 416 360 992 440
rect 416 440 992 520
rect 416 520 992 600
rect 416 600 992 680
rect 416 680 992 760
<< ntap >>
rect -96 -40 96 40
rect 1312 -40 1504 40
rect -96 40 96 120
rect 1312 40 1504 120
rect -96 120 96 200
rect 1312 120 1504 200
rect -96 200 96 280
rect 1312 200 1504 280
rect -96 280 96 360
rect 1312 280 1504 360
rect -96 360 96 440
rect 1312 360 1504 440
rect -96 440 96 520
rect 1312 440 1504 520
rect -96 520 96 600
rect 1312 520 1504 600
rect -96 600 96 680
rect 1312 600 1504 680
rect -96 680 96 760
rect 1312 680 1504 760
rect -96 760 96 840
rect 1312 760 1504 840
<< poly >>
rect 160 146 1248 334
rect 160 466 1248 654
rect 160 -22 1248 22
rect 160 200 224 280
rect 1184 200 1248 280
rect 160 280 224 360
rect 1184 280 1248 360
rect 160 360 224 440
rect 1184 360 1248 440
rect 160 440 224 520
rect 1184 440 1248 520
rect 160 520 224 600
rect 1184 520 1248 600
rect 160 778 1248 822
<< m1 >>
rect 160 360 224 440
rect 288 600 480 680
rect 928 40 1120 120
rect 160 40 224 120
rect 288 40 480 120
rect 928 40 1120 120
rect 160 120 224 200
rect 288 120 480 200
rect 928 120 1120 200
rect 160 200 224 280
rect 288 200 480 280
rect 928 200 1120 280
rect 160 280 224 360
rect 288 280 480 360
rect 928 280 1120 360
rect 160 360 224 440
rect 288 360 480 440
rect 928 360 1120 440
rect 160 440 224 520
rect 288 440 480 520
rect 928 440 1120 520
rect 160 520 224 600
rect 288 520 480 600
rect 928 520 1120 600
rect 160 600 224 680
rect 288 600 480 680
rect 928 600 1120 680
rect 160 680 224 760
rect 288 680 480 760
rect 928 680 1120 760
<< pcontact >>
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 1195 300 1237 320
rect 1195 320 1237 340
rect 1195 340 1237 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 1195 360 1237 380
rect 1195 380 1237 400
rect 1195 400 1237 420
rect 1195 420 1237 440
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 1195 440 1237 460
rect 1195 460 1237 480
rect 1195 480 1237 500
<< locali >>
rect -96 -40 96 40
rect 1312 -40 1504 40
rect -96 40 96 120
rect 288 40 992 120
rect 1312 40 1504 120
rect -96 120 96 200
rect 1312 120 1504 200
rect -96 200 96 280
rect 1312 200 1504 280
rect -96 280 96 360
rect 160 280 224 360
rect 1184 280 1248 360
rect 1312 280 1504 360
rect -96 360 96 440
rect -96 360 96 440
rect 160 360 224 440
rect 416 360 1120 440
rect 1184 360 1248 440
rect 1312 360 1504 440
rect -96 440 96 520
rect 160 440 224 520
rect 1184 440 1248 520
rect 1312 440 1504 520
rect -96 520 96 600
rect 1312 520 1504 600
rect -96 600 96 680
rect 1312 600 1504 680
rect -96 680 96 760
rect 288 680 992 760
rect 1312 680 1504 760
rect -96 760 96 840
rect 1312 760 1504 840
<< ntapc >>
rect -32 200 32 280
rect 1376 200 1440 280
rect -32 280 32 360
rect 1376 280 1440 360
rect -32 360 32 440
rect 1376 360 1440 440
rect -32 440 32 520
rect 1376 440 1440 520
rect -32 520 32 600
rect 1376 520 1440 600
<< pdcontact >>
rect 448 60 480 80
rect 448 80 480 100
rect 480 60 544 80
rect 480 80 544 100
rect 544 60 608 80
rect 544 80 608 100
rect 608 60 672 80
rect 608 80 672 100
rect 672 60 736 80
rect 672 80 736 100
rect 736 60 800 80
rect 736 80 800 100
rect 800 60 864 80
rect 800 80 864 100
rect 864 60 928 80
rect 864 80 928 100
rect 928 60 960 80
rect 928 80 960 100
rect 448 380 480 400
rect 448 400 480 420
rect 480 380 544 400
rect 480 400 544 420
rect 544 380 608 400
rect 544 400 608 420
rect 608 380 672 400
rect 608 400 672 420
rect 672 380 736 400
rect 672 400 736 420
rect 736 380 800 400
rect 736 400 800 420
rect 800 380 864 400
rect 800 400 864 420
rect 864 380 928 400
rect 864 400 928 420
rect 928 380 960 400
rect 928 400 960 420
rect 448 700 480 720
rect 448 720 480 740
rect 480 700 544 720
rect 480 720 544 740
rect 544 700 608 720
rect 544 720 608 740
rect 608 700 672 720
rect 608 720 672 740
rect 672 700 736 720
rect 672 720 736 740
rect 736 700 800 720
rect 736 720 800 740
rect 800 700 864 720
rect 800 720 864 740
rect 864 700 928 720
rect 864 720 928 740
rect 928 700 960 720
rect 928 720 960 740
<< viali >>
rect 320 48 352 56
rect 320 56 352 64
rect 320 64 352 72
rect 320 72 352 80
rect 320 80 352 88
rect 320 88 352 96
rect 320 96 352 104
rect 320 104 352 112
rect 352 48 416 56
rect 352 56 416 64
rect 352 64 416 72
rect 352 72 416 80
rect 352 80 416 88
rect 352 88 416 96
rect 352 96 416 104
rect 352 104 416 112
rect 416 48 448 56
rect 416 56 448 64
rect 416 64 448 72
rect 416 72 448 80
rect 416 80 448 88
rect 416 88 448 96
rect 416 96 448 104
rect 416 104 448 112
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 960 368 992 376
rect 960 376 992 384
rect 960 384 992 392
rect 960 392 992 400
rect 960 400 992 408
rect 960 408 992 416
rect 960 416 992 424
rect 960 424 992 432
rect 992 368 1056 376
rect 992 376 1056 384
rect 992 384 1056 392
rect 992 392 1056 400
rect 992 400 1056 408
rect 992 408 1056 416
rect 992 416 1056 424
rect 992 424 1056 432
rect 1056 368 1088 376
rect 1056 376 1088 384
rect 1056 384 1088 392
rect 1056 392 1088 400
rect 1056 400 1088 408
rect 1056 408 1088 416
rect 1056 416 1088 424
rect 1056 424 1088 432
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 320 688 352 696
rect 320 696 352 704
rect 320 704 352 712
rect 320 712 352 720
rect 320 720 352 728
rect 320 728 352 736
rect 320 736 352 744
rect 320 744 352 752
rect 352 688 416 696
rect 352 696 416 704
rect 352 704 416 712
rect 352 712 416 720
rect 352 720 416 728
rect 352 728 416 736
rect 352 736 416 744
rect 352 744 416 752
rect 416 688 448 696
rect 416 696 448 704
rect 416 704 448 712
rect 416 712 448 720
rect 416 720 448 728
rect 416 728 448 736
rect 416 736 448 744
rect 416 744 448 752
<< pmoslvt >>
rect 416 146 992 334
rect 416 466 992 654
<< nwell >>
rect -184 -128 1592 928
<< labels >>
flabel m1 s 160 360 224 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 288 600 480 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -96 360 96 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 928 40 1120 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -184 -128 1592 928
<< end >>
