magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1336 608
<< ptap >>
rect -96 120 1248 200
rect -96 200 1248 280
rect -96 280 1248 360
rect -96 360 96 440
rect 1056 360 1248 440
rect -96 440 96 520
rect 1056 440 1248 520
<< locali >>
rect -96 120 1248 200
rect -96 200 1248 280
rect -96 280 1248 360
rect -96 360 96 440
rect 1056 360 1248 440
rect -96 440 96 520
rect 1056 440 1248 520
<< ptapc >>
rect 160 200 928 280
<< pwell >>
rect -184 -128 1336 608
<< labels >>
<< properties >>
string FIXED_BBOX -184 -128 1336 608
<< end >>
