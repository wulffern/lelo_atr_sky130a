magic
tech sky130A
magscale 1 2
timestamp 1767481200
<< checkpaint >>
rect -184 -128 1848 928
<< pdiff >>
rect 416 40 1248 120
rect 416 120 1248 200
rect 416 200 1248 280
rect 416 280 1248 360
rect 416 360 1248 440
rect 416 440 1248 520
rect 416 520 1248 600
rect 416 600 1248 680
rect 416 680 1248 760
<< ntap >>
rect -96 -40 96 40
rect 1568 -40 1760 40
rect -96 40 96 120
rect 1568 40 1760 120
rect -96 120 96 200
rect 1568 120 1760 200
rect -96 200 96 280
rect 1568 200 1760 280
rect -96 280 96 360
rect 1568 280 1760 360
rect -96 360 96 440
rect 1568 360 1760 440
rect -96 440 96 520
rect 1568 440 1760 520
rect -96 520 96 600
rect 1568 520 1760 600
rect -96 600 96 680
rect 1568 600 1760 680
rect -96 680 96 760
rect 1568 680 1760 760
rect -96 760 96 840
rect 1568 760 1760 840
<< poly >>
rect 160 146 1504 334
rect 160 466 1504 654
rect 160 -22 1504 22
rect 160 200 224 280
rect 1440 200 1504 280
rect 160 280 224 360
rect 1440 280 1504 360
rect 160 360 224 440
rect 1440 360 1504 440
rect 160 440 224 520
rect 1440 440 1504 520
rect 160 520 224 600
rect 1440 520 1504 600
rect 160 778 1504 822
<< m1 >>
rect 160 360 224 440
rect 288 600 480 680
rect 1184 40 1376 120
rect 160 40 224 120
rect 288 40 480 120
rect 1184 40 1376 120
rect 160 120 224 200
rect 288 120 480 200
rect 1184 120 1376 200
rect 160 200 224 280
rect 288 200 480 280
rect 1184 200 1376 280
rect 160 280 224 360
rect 288 280 480 360
rect 1184 280 1376 360
rect 160 360 224 440
rect 288 360 480 440
rect 1184 360 1376 440
rect 160 440 224 520
rect 288 440 480 520
rect 1184 440 1376 520
rect 160 520 224 600
rect 288 520 480 600
rect 1184 520 1376 600
rect 160 600 224 680
rect 288 600 480 680
rect 1184 600 1376 680
rect 160 680 224 760
rect 288 680 480 760
rect 1184 680 1376 760
<< pcontact >>
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 1451 300 1493 320
rect 1451 320 1493 340
rect 1451 340 1493 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 1451 360 1493 380
rect 1451 380 1493 400
rect 1451 400 1493 420
rect 1451 420 1493 440
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 1451 440 1493 460
rect 1451 460 1493 480
rect 1451 480 1493 500
<< locali >>
rect -96 -40 96 40
rect 1568 -40 1760 40
rect -96 40 96 120
rect 288 40 1248 120
rect 1568 40 1760 120
rect -96 120 96 200
rect 1568 120 1760 200
rect -96 200 96 280
rect 1568 200 1760 280
rect -96 280 96 360
rect 160 280 224 360
rect 1440 280 1504 360
rect 1568 280 1760 360
rect -96 360 96 440
rect -96 360 96 440
rect 160 360 224 440
rect 416 360 1376 440
rect 1440 360 1504 440
rect 1568 360 1760 440
rect -96 440 96 520
rect 160 440 224 520
rect 1440 440 1504 520
rect 1568 440 1760 520
rect -96 520 96 600
rect 1568 520 1760 600
rect -96 600 96 680
rect 1568 600 1760 680
rect -96 680 96 760
rect 288 680 1248 760
rect 1568 680 1760 760
rect -96 760 96 840
rect 1568 760 1760 840
<< ntapc >>
rect -32 200 32 280
rect 1632 200 1696 280
rect -32 280 32 360
rect 1632 280 1696 360
rect -32 360 32 440
rect 1632 360 1696 440
rect -32 440 32 520
rect 1632 440 1696 520
rect -32 520 32 600
rect 1632 520 1696 600
<< pdcontact >>
rect 448 60 480 80
rect 448 80 480 100
rect 480 60 544 80
rect 480 80 544 100
rect 544 60 608 80
rect 544 80 608 100
rect 608 60 672 80
rect 608 80 672 100
rect 672 60 736 80
rect 672 80 736 100
rect 736 60 800 80
rect 736 80 800 100
rect 800 60 864 80
rect 800 80 864 100
rect 864 60 928 80
rect 864 80 928 100
rect 928 60 992 80
rect 928 80 992 100
rect 992 60 1056 80
rect 992 80 1056 100
rect 1056 60 1120 80
rect 1056 80 1120 100
rect 1120 60 1184 80
rect 1120 80 1184 100
rect 1184 60 1216 80
rect 1184 80 1216 100
rect 448 380 480 400
rect 448 400 480 420
rect 480 380 544 400
rect 480 400 544 420
rect 544 380 608 400
rect 544 400 608 420
rect 608 380 672 400
rect 608 400 672 420
rect 672 380 736 400
rect 672 400 736 420
rect 736 380 800 400
rect 736 400 800 420
rect 800 380 864 400
rect 800 400 864 420
rect 864 380 928 400
rect 864 400 928 420
rect 928 380 992 400
rect 928 400 992 420
rect 992 380 1056 400
rect 992 400 1056 420
rect 1056 380 1120 400
rect 1056 400 1120 420
rect 1120 380 1184 400
rect 1120 400 1184 420
rect 1184 380 1216 400
rect 1184 400 1216 420
rect 448 700 480 720
rect 448 720 480 740
rect 480 700 544 720
rect 480 720 544 740
rect 544 700 608 720
rect 544 720 608 740
rect 608 700 672 720
rect 608 720 672 740
rect 672 700 736 720
rect 672 720 736 740
rect 736 700 800 720
rect 736 720 800 740
rect 800 700 864 720
rect 800 720 864 740
rect 864 700 928 720
rect 864 720 928 740
rect 928 700 992 720
rect 928 720 992 740
rect 992 700 1056 720
rect 992 720 1056 740
rect 1056 700 1120 720
rect 1056 720 1120 740
rect 1120 700 1184 720
rect 1120 720 1184 740
rect 1184 700 1216 720
rect 1184 720 1216 740
<< viali >>
rect 320 48 352 56
rect 320 56 352 64
rect 320 64 352 72
rect 320 72 352 80
rect 320 80 352 88
rect 320 88 352 96
rect 320 96 352 104
rect 320 104 352 112
rect 352 48 416 56
rect 352 56 416 64
rect 352 64 416 72
rect 352 72 416 80
rect 352 80 416 88
rect 352 88 416 96
rect 352 96 416 104
rect 352 104 416 112
rect 416 48 448 56
rect 416 56 448 64
rect 416 64 448 72
rect 416 72 448 80
rect 416 80 448 88
rect 416 88 448 96
rect 416 96 448 104
rect 416 104 448 112
rect 171 300 213 320
rect 171 320 213 340
rect 171 340 213 360
rect 171 360 213 380
rect 171 380 213 400
rect 171 400 213 420
rect 171 420 213 440
rect 1216 368 1248 376
rect 1216 376 1248 384
rect 1216 384 1248 392
rect 1216 392 1248 400
rect 1216 400 1248 408
rect 1216 408 1248 416
rect 1216 416 1248 424
rect 1216 424 1248 432
rect 1248 368 1312 376
rect 1248 376 1312 384
rect 1248 384 1312 392
rect 1248 392 1312 400
rect 1248 400 1312 408
rect 1248 408 1312 416
rect 1248 416 1312 424
rect 1248 424 1312 432
rect 1312 368 1344 376
rect 1312 376 1344 384
rect 1312 384 1344 392
rect 1312 392 1344 400
rect 1312 400 1344 408
rect 1312 408 1344 416
rect 1312 416 1344 424
rect 1312 424 1344 432
rect 171 440 213 460
rect 171 460 213 480
rect 171 480 213 500
rect 320 688 352 696
rect 320 696 352 704
rect 320 704 352 712
rect 320 712 352 720
rect 320 720 352 728
rect 320 728 352 736
rect 320 736 352 744
rect 320 744 352 752
rect 352 688 416 696
rect 352 696 416 704
rect 352 704 416 712
rect 352 712 416 720
rect 352 720 416 728
rect 352 728 416 736
rect 352 736 416 744
rect 352 744 416 752
rect 416 688 448 696
rect 416 696 448 704
rect 416 704 448 712
rect 416 712 448 720
rect 416 720 448 728
rect 416 728 448 736
rect 416 736 448 744
rect 416 744 448 752
<< nwell >>
rect -184 -128 1848 928
<< labels >>
flabel m1 s 160 360 224 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 288 600 480 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -96 360 96 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 1184 40 1376 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -184 -128 1848 928
<< end >>
